`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/24/2025 02:30:20 AM
// Design Name: 
// Module Name: ALU_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module ALU_testbench;
wire [15:0] Result;
wire [5:0] Status;
reg [15:0] A,B;
reg [4:0] F;
reg Cin;
ALU_16_bits uut(Result,Status,A,B,F,Cin);
initial begin
    #400 $finish;
end

initial fork 
    //UNUSED OPERATIONS
    #0  {A,B,F,Cin} = {16'hf000,16'h0000,5'b00000,1'b1};
    #10 {A,B,F,Cin} = {16'hf000,16'h0000,5'b00010,1'b1};
    //INC
    #20 {A,B,F,Cin} = {16'h0000,16'h0000,5'b00001,1'b1};
    #30 {A,B,F,Cin} = {16'h0001,16'h0000,5'b00001,1'b1};
    //DEC
    #40 {A,B,F,Cin} = {16'h0001,16'h0000,5'b00011,1'b1};
    //ADD
    #50 {A,B,F,Cin} = {16'h0003,16'h0004,5'b00100,1'b1};
    //ADC
    #60 {A,B,F,Cin} = {16'h0003,16'h0004,5'b00101,1'b1};
    //SUB
    #70 {A,B,F,Cin} = {16'hfffe,16'hffff,5'b00110,1'b1};
    //SBB
    #80 {A,B,F,Cin} = {16'h0007,16'h0003,5'b00111,1'b1};
    //AND
    #90 {A,B,F,Cin} = {16'h0007,16'h0003,5'b01000,1'b1};
    //OR
    #100 {A,B,F,Cin} = {16'h0007,16'h0003,5'b01001,1'b1};
    //XOR
    #110 {A,B,F,Cin} = {16'h0007,16'h0003,5'b01010,1'b1};
    ///NOT
    #120 {A,B,F,Cin} = {16'h0007,16'h0003,5'b01011,1'b1};
    //SHL
    #130 {A,B,F,Cin} = {16'h80f0,16'h0003,5'b10000,1'b1};
    #140 {A,B,F,Cin} = {16'h7521,16'h0003,5'b10000,1'b1};
    //SHR
    #150 {A,B,F,Cin} = {16'h0f0f,16'h0003,5'b10001,1'b1};
    #160 {A,B,F,Cin} = {16'h7521,16'h0003,5'b10001,1'b1};
    //SAL
    #170 {A,B,F,Cin} = {16'hf0f0,16'h0003,5'b10010,1'b1};
    //SAR
    #180 {A,B,F,Cin} = {16'hf0f1,16'h0003,5'b10011,1'b1};
    #190 {A,B,F,Cin} = {16'h7521,16'h0003,5'b10011,1'b1};
    //ROL
    #200 {A,B,F,Cin} = {16'hf0f0,16'h0003,5'b10100,1'b1};
    #210 {A,B,F,Cin} = {16'h7521,16'h0003,5'b10100,1'b1};
    //ROR
    #220 {A,B,F,Cin} = {16'h0f0f,16'h0003,5'b10101,1'b1};
    #230 {A,B,F,Cin} = {16'h7521,16'h0003,5'b10101,1'b1};
    //RCL
    #240 {A,B,F,Cin} = {16'h0f0f,16'h0003,5'b10110,1'b1};
    #250 {A,B,F,Cin} = {16'h7521,16'h0003,5'b10110,1'b1};
    //RCR
    #260 {A,B,F,Cin} = {16'h3f00,16'h0003,5'b10111,1'b1};
    #270 {A,B,F,Cin} = {16'h8f00,16'h0003,5'b10111,1'b1};
    #280 {A,B,F,Cin} = {16'hcf00,16'h0003,5'b10111,1'b1};
    #290 {A,B,F,Cin} = {16'h0f00,16'h0003,5'b10111,1'b1};
    //OVERFLOW FLAG 
    #300 {A,B,F,Cin} = {16'h7ff0,16'h0001,5'b00100,1'b1};
    #310 {A,B,F,Cin} = {16'h7f5f,16'h0001,5'b00101,1'b1};
    #320 {A,B,F,Cin} = {16'h7fcf,16'hfccf,5'b00110,1'b1};
    #330 {A,B,F,Cin} = {16'h7ffb,16'hff45,5'b00111,1'b1};
    //AUX FLAG
    #340 {A,B,F,Cin} = {16'h0004,16'h0005,5'b00110,1'b0};
    #350 {A,B,F,Cin} = {16'h0008,16'h0009,5'b00111,1'b1};
    #360 {A,B,F,Cin} = {16'h0030,16'h0000,5'b00011,1'b0};
    #370 {A,B,F,Cin} = {16'h0009,16'h0008,5'b00100,1'b0};
    #380 {A,B,F,Cin} = {16'h0008,16'h0008,5'b00101,1'b1};
    #390 {A,B,F,Cin} = {16'h000F,16'h0000,5'b00001,1'b0};
join
endmodule